(* keep_hierarchy *)
module top (in1, in2, clk1, clk2, clk3, out);
  input in1, in2, clk1, clk2, clk3;
  output out;
  wire r1q, r2q, u1z, u2z;

  (* keep *) DFF_X1 r1 (.D(in1), .CK(clk1), .Q(r1q));
  (* keep *) DFF_X1 r2 (.D(in2), .CK(clk2), .Q(r2q));
  (* keep *) BUF_X1 u1 (.A(r2q), .Z(u1z));
  (* keep *) AND2_X1 u2 (.A1(r1q), .A2(u1z), .ZN(u2z));
  (* keep *) DFF_X1 r3 (.D(u2z), .CK(clk3), .Q(out));
endmodule
